// assigment_luis1.v
// Temporary top-level wrapper (we will connect real modules later)

module assigment_luis1 (
    input  wire clk,      // placeholder clock
    input  wire reset_n   // placeholder reset (active low)
    // TODO: add switches, keys, HEX, LEDs later
);

    // For now, no internal logic.
    // This is just to satisfy the top-level entity requirement.

endmodule
